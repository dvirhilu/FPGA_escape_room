package constants;

// this package contains references to constants defined by systemverilog localparams
`include "ASCII_chars.svh"
`include "audio_controller_const.svh"

endpackage : constants