package type_definitions;

// package to store user defined SV types
'include "data_transactions.svh"

endpackage : type_definitions