package constants;

// this package contains references to constants defined by systemverilog localparams
`include "ASCII_chars.svh"

endpackage : constants