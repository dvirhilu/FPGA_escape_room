`ifndef ascii_chars
`define ascii_chars
//Character definitions

//numbers
localparam character_0 =8'h30;
localparam character_1 =8'h31;
localparam character_2 =8'h32;
localparam character_3 =8'h33;
localparam character_4 =8'h34;
localparam character_5 =8'h35;
localparam character_6 =8'h36;
localparam character_7 =8'h37;
localparam character_8 =8'h38;
localparam character_9 =8'h39;


//Uppercase Letters
localparam character_A =8'h41;
localparam character_B =8'h42;
localparam character_C =8'h43;
localparam character_D =8'h44;
localparam character_E =8'h45;
localparam character_F =8'h46;
localparam character_G =8'h47;
localparam character_H =8'h48;
localparam character_I =8'h49;
localparam character_J =8'h4A;
localparam character_K =8'h4B;
localparam character_L =8'h4C;
localparam character_M =8'h4D;
localparam character_N =8'h4E;
localparam character_O =8'h4F;
localparam character_P =8'h50;
localparam character_Q =8'h51;
localparam character_R =8'h52;
localparam character_S =8'h53;
localparam character_T =8'h54;
localparam character_U =8'h55;
localparam character_V =8'h56;
localparam character_W =8'h57;
localparam character_X =8'h58;
localparam character_Y =8'h59;
localparam character_Z =8'h5A;

//Lowercase Letters
localparam character_lowercase_a= 8'h61;
localparam character_lowercase_b= 8'h62;
localparam character_lowercase_c= 8'h63;
localparam character_lowercase_d= 8'h64;
localparam character_lowercase_e= 8'h65;
localparam character_lowercase_f= 8'h66;
localparam character_lowercase_g= 8'h67;
localparam character_lowercase_h= 8'h68;
localparam character_lowercase_i= 8'h69;
localparam character_lowercase_j= 8'h6A;
localparam character_lowercase_k= 8'h6B;
localparam character_lowercase_l= 8'h6C;
localparam character_lowercase_m= 8'h6D;
localparam character_lowercase_n= 8'h6E;
localparam character_lowercase_o= 8'h6F;
localparam character_lowercase_p= 8'h70;
localparam character_lowercase_q= 8'h71;
localparam character_lowercase_r= 8'h72;
localparam character_lowercase_s= 8'h73;
localparam character_lowercase_t= 8'h74;
localparam character_lowercase_u= 8'h75;
localparam character_lowercase_v= 8'h76;
localparam character_lowercase_w= 8'h77;
localparam character_lowercase_x= 8'h78;
localparam character_lowercase_y= 8'h79;
localparam character_lowercase_z= 8'h7A;

//Other Characters
localparam character_colon = 8'h3A;          //':'
localparam character_stop = 8'h2E;           //'.'
localparam character_semi_colon = 8'h3B;   //';'
localparam character_minus = 8'h2D;         //'-'
localparam character_divide = 8'h2F;         //'/'
localparam character_plus = 8'h2B;          //'+'
localparam character_comma = 8'h2C;          // ','
localparam character_less_than = 8'h3C;    //'<'
localparam character_greater_than = 8'h3E; //'>'
localparam character_equals = 8'h3D;         //'='
localparam character_question = 8'h3F;      //'?'
localparam character_dollar = 8'h24;         //'$'
localparam character_space=8'h20;           //' '     
localparam character_exclaim=8'h21;          //'!'
`endif